module go_generator(clk,value,data);
input clk;
input [7:0]value;
output reg [15:0]data;
always @(posedge clk)
begin
case (value)
            // Number 1 (G)
	     8'b00010000: data = 16'b0000111111110000;
        8'b00010001: data = 16'b0001111111111000;
        8'b00010010: data = 16'b0011100000011100;
        8'b00010011: data = 16'b0111000000001110;
        8'b00010100: data = 16'b0110000000000110;
        8'b00010101: data = 16'b1110000000000111;
        8'b00010110: data = 16'b1100000000000000;
        8'b00010111: data = 16'b1100000000000000;
        8'b00011000: data = 16'b1100000011111111;
        8'b00011001: data = 16'b1100000011111111;
        8'b00011010: data = 16'b1110000000000111;
        8'b00011011: data = 16'b0110000000000110;
        8'b00011100: data = 16'b0111000000001110;
        8'b00011101: data = 16'b0011100000011100;
        8'b00011110: data = 16'b0001111111111000;
        8'b00011111: data = 16'b0000111111110000;


			// Number 2 (A)
        8'b00100000: data = 16'b0000000111000000;
        8'b00100001: data = 16'b0000001111100000;
        8'b00100010: data = 16'b0000011000110000;
        8'b00100011: data = 16'b0000110000011000;
        8'b00100100: data = 16'b0000110000011000;
        8'b00100101: data = 16'b0001100000001100;
        8'b00100110: data = 16'b0011000000001100;
        8'b00100111: data = 16'b0110000000000110;
        8'b00101000: data = 16'b0110000000000110;
        8'b00101001: data = 16'b1111111111111111;
        8'b00101010: data = 16'b1111111111111111;
        8'b00101011: data = 16'b0110000000000110;
        8'b00101100: data = 16'b0110000000000110;
        8'b00101101: data = 16'b0110000000000110;
        8'b00101110: data = 16'b1111000000001111;
        8'b00101111: data = 16'b1111000000001111;


			// Number 3 (M)
        8'b00110000: data = 16'b1110000000000111;
        8'b00110001: data = 16'b1111000000001111;
        8'b00110010: data = 16'b1111100000011111;
        8'b00110011: data = 16'b1101110000111011;
        8'b00110100: data = 16'b1100111001110011;
        8'b00110101: data = 16'b1100011111100011;
        8'b00110110: data = 16'b1100001111000011;
        8'b00110111: data = 16'b1100000110000011;
        8'b00111000: data = 16'b1100000000000011;
        8'b00111001: data = 16'b1100000000000011;
        8'b00111010: data = 16'b1100000000000011;
        8'b00111011: data = 16'b1100000000000011;
        8'b00111100: data = 16'b1100000000000011;
        8'b00111101: data = 16'b1100000000000011;
        8'b00111110: data = 16'b1100000000000011;
        8'b00111111: data = 16'b1100000000000011;


			// Number 4 (E)
        8'b01000000: data = 16'b1111111111111111;
        8'b01000001: data = 16'b1111111111111111;
        8'b01000010: data = 16'b1100000000000000;
        8'b01000011: data = 16'b1100000000000000;
        8'b01000100: data = 16'b1100000000000000;
        8'b01000101: data = 16'b1100000000000000;
        8'b01000110: data = 16'b1111111111111000;
        8'b01000111: data = 16'b1111111111111000;
        8'b01001000: data = 16'b1100000000000000;
        8'b01001001: data = 16'b1100000000000000;
        8'b01001010: data = 16'b1100000000000000;
        8'b01001011: data = 16'b1100000000000000;
        8'b01001100: data = 16'b1100000000000000;
        8'b01001101: data = 16'b1100000000000000;
        8'b01001110: data = 16'b1111111111111111;
        8'b01001111: data = 16'b1111111111111111;


			// Number 5 (O)
        8'b01010000: data = 16'b0011111111111100;
        8'b01010001: data = 16'b0111111111111110;
        8'b01010010: data = 16'b1110000000000111;
        8'b01010011: data = 16'b1100000000000011;
        8'b01010100: data = 16'b1100000000000011;
        8'b01010101: data = 16'b1100000000000011;
        8'b01010110: data = 16'b1100000000000011;
        8'b01010111: data = 16'b1100000000000011;
        8'b01011000: data = 16'b1100000000000011;
        8'b01011001: data = 16'b1100000000000011;
        8'b01011010: data = 16'b1100000000000011;
        8'b01011011: data = 16'b1100000000000011;
        8'b01011100: data = 16'b1100000000000011;
        8'b01011101: data = 16'b1110000000000111;
        8'b01011110: data = 16'b0111111111111110;
        8'b01011111: data = 16'b0011111111111100;

			
			// Number 6 (V)
        8'b01100000: data = 16'b1100000000000011;
        8'b01100001: data = 16'b1100000000000011;
        8'b01100010: data = 16'b1100000000000011;
        8'b01100011: data = 16'b1100000000000011;
        8'b01100100: data = 16'b1100000000000011;
        8'b01100101: data = 16'b1100000000000011;
        8'b01100110: data = 16'b1100000000000011;
        8'b01100111: data = 16'b1100000000000011;
        8'b01101000: data = 16'b0110000000000110;
        8'b01101001: data = 16'b0110000000000110;
        8'b01101010: data = 16'b0011000000001100;
        8'b01101011: data = 16'b0011000000001100;
        8'b01101100: data = 16'b0001100000011000;
        8'b01101101: data = 16'b0000110000110000;
        8'b01101110: data = 16'b0000011111100000;
        8'b01101111: data = 16'b0000001111000000;


			// Number 7 (R)
        8'b01110000: data = 16'b1111111111111000;
        8'b01110001: data = 16'b1111111111111100;
        8'b01110010: data = 16'b1100000000001110;
        8'b01110011: data = 16'b1100000000000111;
        8'b01110100: data = 16'b1100000000000111;
        8'b01110101: data = 16'b1100000000000111;
        8'b01110110: data = 16'b1100000000001110;
        8'b01110111: data = 16'b1100000000011100;
        8'b01111000: data = 16'b1111111111111000;
        8'b01111001: data = 16'b1111111111100000;
        8'b01111010: data = 16'b1100000011100000;
        8'b01111011: data = 16'b1100000001110000;
        8'b01111100: data = 16'b1100000000111000;
        8'b01111101: data = 16'b1100000000011100;
        8'b01111110: data = 16'b1100000000001110;
        8'b01111111: data = 16'b1100000000000111;


//			// Number 8 (1000)
//			8'b10000000: data = 8'b01111110;
//			8'b10000001: data = 8'b01111110;
//			8'b10000010: data = 8'b00000110;
//			8'b10000011: data = 8'b00001100;
//			8'b10000100: data = 8'b00001100;
//			8'b10000101: data = 8'b00011000;
//			8'b10000110: data = 8'b00011000;
//			8'b10000111: data = 8'b00011000;
//			8'b10001000: data = 8'b00011000;
//			8'b10001001: data = 8'b00011000;
//			8'b10001010: data = 8'b00000000;
//			8'b10001011: data = 8'b00000000;
//			8'b10001100: data = 8'b00000000;
//			8'b10001101: data = 8'b00000000;
//			8'b10001110: data = 8'b00000000;
//			8'b10001111: data = 8'b00000000;

//			// Number 9 (1001)
//			8'b10010000: data = 8'b00111100;
//			8'b10010001: data = 8'b01111110;
//			8'b10010010: data = 8'b01100110;
//			8'b10010011: data = 8'b01100110;
//			8'b10010100: data = 8'b01111110;
//			8'b10010101: data = 8'b00111100;
//			8'b10010110: data = 8'b01100110;
//			8'b10010111: data = 8'b01100110;
//			8'b10011000: data = 8'b01111110;
//			8'b10011001: data = 8'b00111100;
//			8'b10011010: data = 8'b00000000;
//			8'b10011011: data = 8'b00000000;
//			8'b10011100: data = 8'b00000000;
//			8'b10011101: data = 8'b00000000;
//			8'b10011110: data = 8'b00000000;
//			8'b10011111: data = 8'b00000000;

//			// Number 10 (1010)
//			8'b10100000: data = 8'b00111100;
//			8'b10100001: data = 8'b01111110;
//			8'b10100010: data = 8'b01100110;
//			8'b10100011: data = 8'b01100110;
//			8'b10100100: data = 8'b01111110;
//			8'b10100101: data = 8'b00111110;
//			8'b10100110: data = 8'b00000110;
//			8'b10100111: data = 8'b00000110;
//			8'b10101000: data = 8'b01111110;
//			8'b10101001: data = 8'b00111100;
//			8'b10101010: data = 8'b00000000;
//			8'b10101011: data = 8'b00000000; 
 
            default:data=0;
  
endcase
end
endmodule
